
let max(a,b) = (a > b) ? a : b;
let max3(a,b,c) = (a>b) ? max(a,c) : max(b,c);