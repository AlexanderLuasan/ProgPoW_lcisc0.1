package EV_enums;




typedef enum{
	shared,
	thread,
	data
} register_select_t;






endpackage;
